module hex7seg(SW,HEX);

	input [3:0] SW;
	output [6:0] HEX;
	
	always @*
		case (SW)
		
			4'b0000 : HEX = 7'b0000001;
			4'b0001 : HEX = 7'b1001111;
			4'b0010 : HEX = 7'b0010010; 
			4'b0011 : HEX = 7'b0000110;
			4'b0100 : HEX = 7'b1001100;
			4'b0101 : HEX = 7'b0100100;  
			4'b0110 : HEX = 7'b0100000;
			4'b0111 : HEX = 7'b0001111;
			4'b1000 : HEX = 7'b0000000;
			4'b1001 : HEX = 7'b0000100;
			4'b1010 : HEX = 7'b0001000; 
			4'b1011 : HEX = 7'b1100000;
			4'b1100 : HEX = 7'b0110001;
			4'b1101 : HEX = 7'b1000010;
			4'b1110 : HEX = 7'b0110000;
			4'b1111 : HEX = 7'b0111000;
			
		endcase
			
	
endmodule

